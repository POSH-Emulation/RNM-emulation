../simulation_src/eg.sv